module uut_always01(input in, output out);

assign out = ~in;

endmodule
